module bitwise_or(output[31:0] res, input[31:0] A, input[31:0] B);
    or or0(res[0], A[0], B[0]);
    or or1(res[1], A[1], B[1]);
    or or2(res[2], A[2], B[2]);
    or or3(res[3], A[3], B[3]);
    or or4(res[4], A[4], B[4]);
    or or5(res[5], A[5], B[5]);
    or or6(res[6], A[6], B[6]);
    or or7(res[7], A[7], B[7]);
    or or8(res[8], A[8], B[8]);
    or or9(res[9], A[9], B[9]);
    or or10(res[10], A[10], B[10]);
    or or11(res[11], A[11], B[11]);
    or or12(res[12], A[12], B[12]);
    or or13(res[13], A[13], B[13]);
    or or14(res[14], A[14], B[14]);
    or or15(res[15], A[15], B[15]);
    or or16(res[16], A[16], B[16]);
    or or17(res[17], A[17], B[17]);
    or or18(res[18], A[18], B[18]);
    or or19(res[19], A[19], B[19]);
    or or20(res[20], A[20], B[20]);
    or or21(res[21], A[21], B[21]);
    or or22(res[22], A[22], B[22]);
    or or23(res[23], A[23], B[23]);
    or or24(res[24], A[24], B[24]);
    or or25(res[25], A[25], B[25]);
    or or26(res[26], A[26], B[26]);
    or or27(res[27], A[27], B[27]);
    or or28(res[28], A[28], B[28]);
    or or29(res[29], A[29], B[29]);
    or or30(res[30], A[30], B[30]);
    or or31(res[31], A[31], B[31]);
endmodule