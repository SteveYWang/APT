module multException(
    output exception,
    input[64:0] finalProd,
    input signA, signB
);
    wire isOne, isZero, sign, isMaxNeg, sameSign;
    assign sign = finalProd[32];
    assign sameSign = (signA & signB) | (~signA & ~signB);

    or or1(isOne,
        finalProd[62],
        finalProd[61],
        finalProd[60],
        finalProd[59],
        finalProd[58],
        finalProd[57],
        finalProd[56],
        finalProd[55],
        finalProd[54],
        finalProd[53],
        finalProd[52],
        finalProd[51],
        finalProd[50],
        finalProd[49],
        finalProd[48],
        finalProd[47],
        finalProd[46],
        finalProd[45],
        finalProd[44],
        finalProd[43],
        finalProd[42],
        finalProd[41],
        finalProd[40],
        finalProd[39],
        finalProd[38],
        finalProd[37],
        finalProd[36],
        finalProd[35],
        finalProd[34],
        finalProd[33]
        );

    or or2(isZero,
        ~finalProd[62],  
        ~finalProd[61],  
        ~finalProd[60],  
        ~finalProd[59],  
        ~finalProd[58],  
        ~finalProd[57],  
        ~finalProd[56],  
        ~finalProd[55],  
        ~finalProd[54],  
        ~finalProd[53],  
        ~finalProd[52],  
        ~finalProd[51],  
        ~finalProd[50],  
        ~finalProd[49],  
        ~finalProd[48],  
        ~finalProd[47],  
        ~finalProd[46],  
        ~finalProd[45],  
        ~finalProd[44],  
        ~finalProd[43],  
        ~finalProd[42],  
        ~finalProd[41],  
        ~finalProd[40],  
        ~finalProd[39],  
        ~finalProd[38],  
        ~finalProd[37],  
        ~finalProd[36],  
        ~finalProd[35],  
        ~finalProd[34],  
        ~finalProd[33]
        );

    and and1(isMaxNeg,
            finalProd[32],
            ~finalProd[31],
            ~finalProd[30],
            ~finalProd[29],
            ~finalProd[28],
            ~finalProd[27],
            ~finalProd[26],
            ~finalProd[25],
            ~finalProd[24],
            ~finalProd[23],
            ~finalProd[22],
            ~finalProd[21],
            ~finalProd[20],
            ~finalProd[19],
            ~finalProd[18],
            ~finalProd[17],
            ~finalProd[16],
            ~finalProd[15],
            ~finalProd[14],
            ~finalProd[13],
            ~finalProd[12],
            ~finalProd[11],
            ~finalProd[10],
            ~finalProd[9],
            ~finalProd[8],
            ~finalProd[7],
            ~finalProd[6],
            ~finalProd[5],
            ~finalProd[4],
            ~finalProd[3],
            ~finalProd[2],
            ~finalProd[1]
        );


    assign exception = (~isMaxNeg & ((isOne & ~sign) | (isZero & sign))) | (isMaxNeg & sameSign) ;

endmodule