module isEqual(output out, input[31:0] A, input[31:0] B);
    assign out = ~(A[31] ^ B[31]) &
                ~(A[30] ^ B[30]) &
                ~(A[29] ^ B[29]) &
                ~(A[28] ^ B[28]) &
                ~(A[27] ^ B[27]) &
                ~(A[26] ^ B[26]) &
                ~(A[25] ^ B[25]) &
                ~(A[24] ^ B[24]) &
                ~(A[23] ^ B[23]) &
                ~(A[22] ^ B[22]) &
                ~(A[21] ^ B[21]) &
                ~(A[20] ^ B[20]) &
                ~(A[19] ^ B[19]) &
                ~(A[18] ^ B[18]) &
                ~(A[17] ^ B[17]) &
                ~(A[16] ^ B[16]) &
                ~(A[15] ^ B[15]) &
                ~(A[14] ^ B[14]) &
                ~(A[13] ^ B[13]) &
                ~(A[12] ^ B[12]) &
                ~(A[11] ^ B[11]) &
                ~(A[10] ^ B[10]) &
                ~(A[9] ^ B[9]) &
                ~(A[8] ^ B[8]) &
                ~(A[7] ^ B[7]) &
                ~(A[6] ^ B[6]) &
                ~(A[5] ^ B[5]) &
                ~(A[4] ^ B[4]) &
                ~(A[3] ^ B[3]) &
                ~(A[2] ^ B[2]) &
                ~(A[1] ^ B[1]) &
                ~(A[0] ^ B[0]);
endmodule
