module bitwise_invert(output[31:0] res, input[31:0] A);
    invert invert0(res[0], A[0]);
    invert invert1(res[1], A[1]);
    invert invert2(res[2], A[2]);
    invert invert3(res[3], A[3]);
    invert invert4(res[4], A[4]);
    invert invert5(res[5], A[5]);
    invert invert6(res[6], A[6]);
    invert invert7(res[7], A[7]);
    invert invert8(res[8], A[8]);
    invert invert9(res[9], A[9]);
    invert invert10(res[10], A[10]);
    invert invert11(res[11], A[11]);
    invert invert12(res[12], A[12]);
    invert invert13(res[13], A[13]);
    invert invert14(res[14], A[14]);
    invert invert15(res[15], A[15]);
    invert invert16(res[16], A[16]);
    invert invert17(res[17], A[17]);
    invert invert18(res[18], A[18]);
    invert invert19(res[19], A[19]);
    invert invert20(res[20], A[20]);
    invert invert21(res[21], A[21]);
    invert invert22(res[22], A[22]);
    invert invert23(res[23], A[23]);
    invert invert24(res[24], A[24]);
    invert invert25(res[25], A[25]);
    invert invert26(res[26], A[26]);
    invert invert27(res[27], A[27]);
    invert invert28(res[28], A[28]);
    invert invert29(res[29], A[29]);
    invert invert30(res[30], A[30]);
    invert invert31(res[31], A[31]);
endmodule