module bitwise_and(output[31:0] res, input[31:0] A, input[31:0] B);
    and and0(res[0], A[0], B[0]);
    and and1(res[1], A[1], B[1]);
    and and2(res[2], A[2], B[2]);
    and and3(res[3], A[3], B[3]);
    and and4(res[4], A[4], B[4]);
    and and5(res[5], A[5], B[5]);
    and and6(res[6], A[6], B[6]);
    and and7(res[7], A[7], B[7]);
    and and8(res[8], A[8], B[8]);
    and and9(res[9], A[9], B[9]);
    and and10(res[10], A[10], B[10]);
    and and11(res[11], A[11], B[11]);
    and and12(res[12], A[12], B[12]);
    and and13(res[13], A[13], B[13]);
    and and14(res[14], A[14], B[14]);
    and and15(res[15], A[15], B[15]);
    and and16(res[16], A[16], B[16]);
    and and17(res[17], A[17], B[17]);
    and and18(res[18], A[18], B[18]);
    and and19(res[19], A[19], B[19]);
    and and20(res[20], A[20], B[20]);
    and and21(res[21], A[21], B[21]);
    and and22(res[22], A[22], B[22]);
    and and23(res[23], A[23], B[23]);
    and and24(res[24], A[24], B[24]);
    and and25(res[25], A[25], B[25]);
    and and26(res[26], A[26], B[26]);
    and and27(res[27], A[27], B[27]);
    and and28(res[28], A[28], B[28]);
    and and29(res[29], A[29], B[29]);
    and and30(res[30], A[30], B[30]);
    and and31(res[31], A[31], B[31]);
endmodule